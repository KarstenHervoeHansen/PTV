--
-- VROM initialization values for synthesis
-- Created from file PAL_EG1_RP178.txt on Fri 27 Aug 2004 14:54
-- Formatted for Xilinx XST synthesis tool.
--
attribute WRITE_MODE_A of VROM : label is "READ_FIRST";
attribute WRITE_MODE_B of VROM : label is "READ_FIRST";
attribute INIT_A of VROM : label is "30671";
attribute INIT_B of VROM : label is "30671";
attribute SRVAL_A of VROM : label is "30671";
attribute SRVAL_B of VROM : label is "30671";
attribute INITP_00 of VROM : label is "0000000000000000000000000000000000000000000000000000055555555557";
attribute INITP_01 of VROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_02 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAABFFFFFFFFFFF5000000000000000000000000000";
attribute INITP_03 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_04 of VROM : label is "FFFFFFF7EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_05 of VROM : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
attribute INITP_06 of VROM : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
attribute INITP_07 of VROM : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
attribute INIT_00 of VROM : label is "0010000F000E000D000C000B000A000900080007000600050004000300020671";
attribute INIT_01 of VROM : label is "0C200C1F0C1E0C1D0C1C0C1B0C1A0C190C180817001600150014001300120011";
attribute INIT_02 of VROM : label is "0C300C2F0C2E0C2D0C2C0C2B0C2A0C290C280C270C260C250C240C230C220C21";
attribute INIT_03 of VROM : label is "0C400C3F0C3E0C3D0C3C0C3B0C3A0C390C380C370C360C350C340C330C320C31";
attribute INIT_04 of VROM : label is "0C500C4F0C4E0C4D0C4C0C4B0C4A0C490C480C470C460C450C440C430C420C41";
attribute INIT_05 of VROM : label is "0C600C5F0C5E0C5D0C5C0C5B0C5A0C590C580C570C560C550C540C530C520C51";
attribute INIT_06 of VROM : label is "0C700C6F0C6E0C6D0C6C0C6B0C6A0C690C680C670C660C650C640C630C620C61";
attribute INIT_07 of VROM : label is "0C800C7F0C7E0C7D0C7C0C7B0C7A0C790C780C770C760C750C740C730C720C71";
attribute INIT_08 of VROM : label is "0C900C8F0C8E0C8D0C8C0C8B0C8A0C890C880C870C860C850C840C830C820C81";
attribute INIT_09 of VROM : label is "0CA00C9F0C9E0C9D0C9C0C9B0C9A0C990C980C970C960C950C940C930C920C91";
attribute INIT_0A of VROM : label is "10B010AF10AE10AD10AC10AB10AA10A910A810A710A610A510A410A310A210A1";
attribute INIT_0B of VROM : label is "10C010BF10BE10BD10BC10BB10BA10B910B810B710B610B510B410B310B210B1";
attribute INIT_0C of VROM : label is "10D010CF10CE10CD10CC10CB10CA10C910C810C710C610C510C410C310C210C1";
attribute INIT_0D of VROM : label is "14E014DF14DE14DD14DC14DB14DA14D914D810D710D610D510D410D310D210D1";
attribute INIT_0E of VROM : label is "18F018EF14EE14ED14EC14EB14EA14E914E814E714E614E514E414E314E214E1";
attribute INIT_0F of VROM : label is "190018FF18FE18FD18FC18FB18FA18F918F818F718F618F518F418F318F218F1";
attribute INIT_10 of VROM : label is "1910190F190E190D190C190B190A190919081907190619051904190319021901";
attribute INIT_11 of VROM : label is "1920191F191E191D191C191B191A191919181917191619151914191319121911";
attribute INIT_12 of VROM : label is "1930192F192E192D192C192B192A192919281927192619251924192319221921";
attribute INIT_13 of VROM : label is "0540053F053E053D053C053B053A053901380137193619351934193319321931";
attribute INIT_14 of VROM : label is "1D50054F054E054D054C054B054A054905480547054605450544054305420541";
attribute INIT_15 of VROM : label is "1D601D5F1D5E1D5D1D5C1D5B1D5A1D591D581D571D561D551D541D531D521D51";
attribute INIT_16 of VROM : label is "1D701D6F1D6E1D6D1D6C1D6B1D6A1D691D681D671D661D651D641D631D621D61";
attribute INIT_17 of VROM : label is "1D801D7F1D7E1D7D1D7C1D7B1D7A1D791D781D771D761D751D741D731D721D71";
attribute INIT_18 of VROM : label is "1D901D8F1D8E1D8D1D8C1D8B1D8A1D891D881D871D861D851D841D831D821D81";
attribute INIT_19 of VROM : label is "1DA01D9F1D9E1D9D1D9C1D9B1D9A1D991D981D971D961D951D941D931D921D91";
attribute INIT_1A of VROM : label is "1DB01DAF1DAE1DAD1DAC1DAB1DAA1DA91DA81DA71DA61DA51DA41DA31DA21DA1";
attribute INIT_1B of VROM : label is "1DC01DBF1DBE1DBD1DBC1DBB1DBA1DB91DB81DB71DB61DB51DB41DB31DB21DB1";
attribute INIT_1C of VROM : label is "1DD01DCF1DCE1DCD1DCC1DCB1DCA1DC91DC81DC71DC61DC51DC41DC31DC21DC1";
attribute INIT_1D of VROM : label is "21E021DF21DE21DD21DC21DB21DA1DD91DD81DD71DD61DD51DD41DD31DD21DD1";
attribute INIT_1E of VROM : label is "21F021EF21EE21ED21EC21EB21EA21E921E821E721E621E521E421E321E221E1";
attribute INIT_1F of VROM : label is "220021FF21FE21FD21FC21FB21FA21F921F821F721F621F521F421F321F221F1";
attribute INIT_20 of VROM : label is "2210220F220E220D220C220B220A220922082207220622052204220322022201";
attribute INIT_21 of VROM : label is "2620261F261E261D261C261B261A261926182617261626152614261326122611";
attribute INIT_22 of VROM : label is "2A302A2F2A2E2A2D2A2C2A2B2A2A2A292A282627262626252624262326222621";
attribute INIT_23 of VROM : label is "2A402A3F2A3E2A3D2A3C2A3B2A3A2A392A382A372A362A352A342A332A322A31";
attribute INIT_24 of VROM : label is "2A502A4F2A4E2A4D2A4C2A4B2A4A2A492A482A472A462A452A442A432A422A41";
attribute INIT_25 of VROM : label is "2A602A5F2A5E2A5D2A5C2A5B2A5A2A592A582A572A562A552A542A532A522A51";
attribute INIT_26 of VROM : label is "06702A6F2A6E2A6D2A6C2A6B2A6A2A692A682A672A662A652A642A632A622A61";
attribute INIT_27 of VROM : label is "0671067106710671067106710671067106710671067106710671067100010671";
attribute INIT_28 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_29 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_2A of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_2B of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_2C of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_2D of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_2E of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_2F of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_30 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_31 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_32 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_33 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_34 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_35 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_36 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_37 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_38 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_39 of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_3A of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_3B of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_3C of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_3D of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_3E of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
attribute INIT_3F of VROM : label is "0671067106710671067106710671067106710671067106710671067106710671";
