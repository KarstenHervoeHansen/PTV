LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE sinu_data IS
	type sintable is array(0 to 47) of std_logic_vector(23 downto 0);
	type sintable2 is array(0 to 7) of std_logic_vector(23 downto 0);
	
	constant sinu_1k: sintable :=
		("000000000000000000000000",
		"000010000101101010001010",
		"000100001001000001111110",
		"000110000111110111100010",
		"001000000000000000000000",
		"001001101111010111110010",
		"001011010100000100111100",
		"001100101100011001001101",
		"001101110110110011110101",
		"001110110010000011010111",
		"001111011101000110111010",
		"001111110111001111010101",
		"010000000000000000000000",
		"001111110111001111010101",
		"001111011101000110111010",
		"001110110010000011010111",
		"001101110110110011110101",
		"001100101100011001001101",
		"001011010100000100111100",
		"001001101111010111110010",
		"001000000000000000000000",
		"000110000111110111100010",
		"000100001001000001111110",
		"000010000101101010001010",
		"000000000000000000000000",
		"111101111010010101110110",
		"111011110110111110000010",
		"111001111000001000011110",
		"111000000000000000000000",
		"110110010000101000001110",
		"110100101011111011000100",
		"110011010011100110110011",
		"110010001001001100001011",
		"110001001101111100101001",
		"110000100010111001000110",
		"110000001000110000101011",
		"110000000000000000000000",
		"110000001000110000101011",
		"110000100010111001000110",
		"110001001101111100101001",
		"110010001001001100001011",
		"110011010011100110110011",
		"110100101011111011000100",
		"110110010000101000001110",
		"111000000000000000000000",
		"111001111000001000011110",
		"111011110110111110000010",
		"111101111010010101110110");

--constant sinu6k : sintable2 :=
--	("000000000000000000000000",
--     "001011010111000010100011",	 
--	 "001111111111111111111111",
--     "001011010111000010100011",
--	 "000000000000000000000000",
--     "110100101000111101011100",
--	 "110000000000000000000000",
--     "110100101000111101011100",
--	 "111000000000000000000000");
--
--
--
--constant square: sintable2 := 
-- 	(
-- 	 "001111111111111111111111",
-- 	 "001111111111111111111111", 
-- 	 "001111111111111111111111",
-- 	 "001111111111111111111111", 
-- 	 "110000000000000000000000",
-- 	 "110000000000000000000000",
-- 	 "110000000000000000000000",
-- 	 "110000000000000000000000"�
-- 	 );	 

END sinu_data;
PACKAGE BODY sinu_data IS

END sinu_data;

