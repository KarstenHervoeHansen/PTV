		--
		-- Initialize VROM for simulation
		-- Created from file PAL_EG1_RP178.txt on Fri 27 Aug 2004 14:54
		-- Number of patterns = 2, number of hregion bits = 4, number of vregion bits = 4
		--
-- translate_off
		generic map (
			WRITE_MODE_A => "READ_FIRST",
			WRITE_MODE_B => "READ_FIRST",
			INIT_A       => X"30671",
			INIT_B       => X"30671",
			SRVAL_A      => X"30671",
			SRVAL_B      => X"30671",
			INITP_00 => X"0000000000000000000000000000000000000000000000000000055555555557",
			INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_02 => X"AAAAAAAAAAAAAAAAAAAAAAAABFFFFFFFFFFF5000000000000000000000000000",
			INITP_03 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_04 => X"FFFFFFF7EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_05 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
			INITP_06 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
			INITP_07 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
			INIT_00 => X"0010000F000E000D000C000B000A000900080007000600050004000300020671",
			INIT_01 => X"0C200C1F0C1E0C1D0C1C0C1B0C1A0C190C180817001600150014001300120011",
			INIT_02 => X"0C300C2F0C2E0C2D0C2C0C2B0C2A0C290C280C270C260C250C240C230C220C21",
			INIT_03 => X"0C400C3F0C3E0C3D0C3C0C3B0C3A0C390C380C370C360C350C340C330C320C31",
			INIT_04 => X"0C500C4F0C4E0C4D0C4C0C4B0C4A0C490C480C470C460C450C440C430C420C41",
			INIT_05 => X"0C600C5F0C5E0C5D0C5C0C5B0C5A0C590C580C570C560C550C540C530C520C51",
			INIT_06 => X"0C700C6F0C6E0C6D0C6C0C6B0C6A0C690C680C670C660C650C640C630C620C61",
			INIT_07 => X"0C800C7F0C7E0C7D0C7C0C7B0C7A0C790C780C770C760C750C740C730C720C71",
			INIT_08 => X"0C900C8F0C8E0C8D0C8C0C8B0C8A0C890C880C870C860C850C840C830C820C81",
			INIT_09 => X"0CA00C9F0C9E0C9D0C9C0C9B0C9A0C990C980C970C960C950C940C930C920C91",
			INIT_0A => X"10B010AF10AE10AD10AC10AB10AA10A910A810A710A610A510A410A310A210A1",
			INIT_0B => X"10C010BF10BE10BD10BC10BB10BA10B910B810B710B610B510B410B310B210B1",
			INIT_0C => X"10D010CF10CE10CD10CC10CB10CA10C910C810C710C610C510C410C310C210C1",
			INIT_0D => X"14E014DF14DE14DD14DC14DB14DA14D914D810D710D610D510D410D310D210D1",
			INIT_0E => X"18F018EF14EE14ED14EC14EB14EA14E914E814E714E614E514E414E314E214E1",
			INIT_0F => X"190018FF18FE18FD18FC18FB18FA18F918F818F718F618F518F418F318F218F1",
			INIT_10 => X"1910190F190E190D190C190B190A190919081907190619051904190319021901",
			INIT_11 => X"1920191F191E191D191C191B191A191919181917191619151914191319121911",
			INIT_12 => X"1930192F192E192D192C192B192A192919281927192619251924192319221921",
			INIT_13 => X"0540053F053E053D053C053B053A053901380137193619351934193319321931",
			INIT_14 => X"1D50054F054E054D054C054B054A054905480547054605450544054305420541",
			INIT_15 => X"1D601D5F1D5E1D5D1D5C1D5B1D5A1D591D581D571D561D551D541D531D521D51",
			INIT_16 => X"1D701D6F1D6E1D6D1D6C1D6B1D6A1D691D681D671D661D651D641D631D621D61",
			INIT_17 => X"1D801D7F1D7E1D7D1D7C1D7B1D7A1D791D781D771D761D751D741D731D721D71",
			INIT_18 => X"1D901D8F1D8E1D8D1D8C1D8B1D8A1D891D881D871D861D851D841D831D821D81",
			INIT_19 => X"1DA01D9F1D9E1D9D1D9C1D9B1D9A1D991D981D971D961D951D941D931D921D91",
			INIT_1A => X"1DB01DAF1DAE1DAD1DAC1DAB1DAA1DA91DA81DA71DA61DA51DA41DA31DA21DA1",
			INIT_1B => X"1DC01DBF1DBE1DBD1DBC1DBB1DBA1DB91DB81DB71DB61DB51DB41DB31DB21DB1",
			INIT_1C => X"1DD01DCF1DCE1DCD1DCC1DCB1DCA1DC91DC81DC71DC61DC51DC41DC31DC21DC1",
			INIT_1D => X"21E021DF21DE21DD21DC21DB21DA1DD91DD81DD71DD61DD51DD41DD31DD21DD1",
			INIT_1E => X"21F021EF21EE21ED21EC21EB21EA21E921E821E721E621E521E421E321E221E1",
			INIT_1F => X"220021FF21FE21FD21FC21FB21FA21F921F821F721F621F521F421F321F221F1",
			INIT_20 => X"2210220F220E220D220C220B220A220922082207220622052204220322022201",
			INIT_21 => X"2620261F261E261D261C261B261A261926182617261626152614261326122611",
			INIT_22 => X"2A302A2F2A2E2A2D2A2C2A2B2A2A2A292A282627262626252624262326222621",
			INIT_23 => X"2A402A3F2A3E2A3D2A3C2A3B2A3A2A392A382A372A362A352A342A332A322A31",
			INIT_24 => X"2A502A4F2A4E2A4D2A4C2A4B2A4A2A492A482A472A462A452A442A432A422A41",
			INIT_25 => X"2A602A5F2A5E2A5D2A5C2A5B2A5A2A592A582A572A562A552A542A532A522A51",
			INIT_26 => X"06702A6F2A6E2A6D2A6C2A6B2A6A2A692A682A672A662A652A642A632A622A61",
			INIT_27 => X"0671067106710671067106710671067106710671067106710671067100010671",
			INIT_28 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_29 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_2A => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_2B => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_2C => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_2D => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_2E => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_2F => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_30 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_31 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_32 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_33 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_34 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_35 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_36 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_37 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_38 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_39 => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_3A => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_3B => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_3C => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_3D => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_3E => X"0671067106710671067106710671067106710671067106710671067106710671",
			INIT_3F => X"0671067106710671067106710671067106710671067106710671067106710671"
		)
-- translate_on
