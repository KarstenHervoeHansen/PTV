--
-- CROM initialization values for synthesis
-- Created from file NTSC_EG1_RP178.txt on Wed 28 Nov 2001 16:12
-- Formatted for Xilinx XST synthesis tool.
--
attribute WRITE_MODE_A of CROM : label is "READ_FIRST";
attribute WRITE_MODE_B of CROM : label is "READ_FIRST";
attribute INIT_A of CROM : label is "000";
attribute INIT_B of CROM : label is "000";
attribute SRVAL_A of CROM : label is "000";
attribute SRVAL_B of CROM : label is "000";
attribute INITP_00 of CROM : label is "995114445AABBEEF995114445AABBEEF99555555555555559955555555555555";
attribute INITP_01 of CROM : label is "9955555555555555995555555555FF11995FF555B5555551995114445AABBEEF";
attribute INITP_02 of CROM : label is "995FF555B5555551995114445AABBEEF995114445AABBEEF9955555555555555";
attribute INITP_03 of CROM : label is "000000000000000000000000000000000000000000000000995555555555FF11";
attribute INITP_04 of CROM : label is "9955555555555555995555555555555599555555555555559955555555555555";
attribute INITP_05 of CROM : label is "9955555555555555995555555555555599555555555555559955555555555555";
attribute INITP_06 of CROM : label is "9955555555555555995555555555555599555555555555559955555555555555";
attribute INITP_07 of CROM : label is "0000000000000000000000000000000000000000000000009955555555555555";
attribute INIT_00 of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_01 of CROM : label is "D80000FFE20000FF200020002000200020002000200020002000200020002000";
attribute INIT_02 of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_03 of CROM : label is "560000FF6C0000FF200020002000200020002000200020002000200020002000";
attribute INIT_04 of CROM : label is "7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800";
attribute INIT_05 of CROM : label is "000000FF3A0000FF2000200037F037A837F037A866A866D966A866D966A866D9";
attribute INIT_06 of CROM : label is "7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800";
attribute INIT_07 of CROM : label is "000000FF3A0000FF2000200037F037A837F037A866A866D966A866D966A866D9";
attribute INIT_08 of CROM : label is "7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800";
attribute INIT_09 of CROM : label is "000000FF3A0000FF2000200037F037A837F037A866A866D966A866D966A866D9";
attribute INIT_0A of CROM : label is "2258222620002000200020007D987D817D987D81200020002000200037F037A8";
attribute INIT_0B of CROM : label is "000000FF3A0000FF200020006800680068006800200020002000200020002000";
attribute INIT_0C of CROM : label is "2000200020002000462F465C462F465CD600D600D600D6007AC57A327AC57A32";
attribute INIT_0D of CROM : label is "000000FF3A0000FF20002000200020002000200031003100200020000E000E00";
attribute INIT_0E of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_0F of CROM : label is "560000FF6C0000FF200020002000200020002000200020002000200020002000";
attribute INIT_10 of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_11 of CROM : label is "D80000FFE20000FF200020002000200020002000200020002000200020002000";
attribute INIT_12 of CROM : label is "7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800";
attribute INIT_13 of CROM : label is "8E0000FFB40000FF2000200037F037A837F037A866A866D966A866D966A866D9";
attribute INIT_14 of CROM : label is "7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800";
attribute INIT_15 of CROM : label is "8E0000FFB40000FF2000200037F037A837F037A866A866D966A866D966A866D9";
attribute INIT_16 of CROM : label is "2258222620002000200020007D987D817D987D81200020002000200037F037A8";
attribute INIT_17 of CROM : label is "8E0000FFB40000FF200020006800680068006800200020002000200020002000";
attribute INIT_18 of CROM : label is "2000200020002000462F465C462F465CD600D600D600D6007AC57A327AC57A32";
attribute INIT_19 of CROM : label is "8E0000FFB40000FF20002000200020002000200031003100200020000E000E00";
attribute INIT_1A of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_21 of CROM : label is "D80000FFE20000FF200020002000200020002000200020002000200020002000";
attribute INIT_22 of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_23 of CROM : label is "560000FF6C0000FF200020002000200020002000200020002000200020002000";
attribute INIT_24 of CROM : label is "CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80";
attribute INIT_25 of CROM : label is "000000FF3A0000FF200020004080CC80CC80CC80CC80CC80CC80CC80CC80CC80";
attribute INIT_26 of CROM : label is "CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80";
attribute INIT_27 of CROM : label is "000000FF3A0000FF20002000CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80";
attribute INIT_28 of CROM : label is "8800880088008800880088008800880088008800880088008800880088008800";
attribute INIT_29 of CROM : label is "000000FF3A0000FF200020008800880088008800880088008800880088008800";
attribute INIT_2A of CROM : label is "8800880088008800880088008800880088008800880088008800880088008800";
attribute INIT_2B of CROM : label is "000000FF3A0000FF200020008800880088008800880088008800880088008800";
attribute INIT_2C of CROM : label is "8800880088008800880088008800880088008800880088008800880088008800";
attribute INIT_2D of CROM : label is "000000FF3A0000FF200020008800880088008800880088008800880088008800";
attribute INIT_2E of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_2F of CROM : label is "560000FF6C0000FF200020002000200020002000200020002000200020002000";
attribute INIT_30 of CROM : label is "2000200020002000200020002000200020002000200020002000200020002000";
attribute INIT_31 of CROM : label is "D80000FFE20000FF200020002000200020002000200020002000200020002000";
attribute INIT_32 of CROM : label is "CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80";
attribute INIT_33 of CROM : label is "8E0000FFB40000FF20002000CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80";
attribute INIT_34 of CROM : label is "8800880088008800880088008800880088008800880088008800880088008800";
attribute INIT_35 of CROM : label is "8E0000FFB40000FF200020008800880088008800880088008800880088008800";
attribute INIT_36 of CROM : label is "8800880088008800880088008800880088008800880088008800880088008800";
attribute INIT_37 of CROM : label is "8E0000FFB40000FF200020008800880088008800880088008800880088008800";
attribute INIT_38 of CROM : label is "8800880088008800880088008800880088008800880088008800880088008800";
attribute INIT_39 of CROM : label is "8E0000FFB40000FF200020008800880088008800880088008800880088008800";
attribute INIT_3A of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of CROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
