		--
		-- Initialize HROM for simulation
		-- Created from file NTSC_EG1_RP178.txt on Wed 28 Nov 2001 16:12
		-- Number of patterns = 2, number of hregion bits = 4, number of vregion bits = 4
		--
-- translate_off
		generic map (
			WRITE_MODE_A => "READ_FIRST",
			WRITE_MODE_B => "READ_FIRST",
			INIT_A       => X"23167",
			INIT_B       => X"23167",
			SRVAL_A      => X"23167",
			SRVAL_B      => X"23167",
			INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_02 => X"5555555555556000000000000000000000000000000000000000000000000000",
			INITP_03 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA85555555555555555555555",
			INITP_04 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_05 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_06 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_07 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INIT_00 => X"0010000F000E000D000C000B000A000900080007000600050004000300020001",
			INIT_01 => X"0020001F001E001D001C001B001A001900180017001600150014001300120011",
			INIT_02 => X"0030002F002E002D002C002B002A002900280027002600250024002300220021",
			INIT_03 => X"0440043F043E043D043C043B043A043904380437043604350434003300320031",
			INIT_04 => X"0850084F084E084D084C084B084A084908480847084608450844084308420841",
			INIT_05 => X"0860085F085E085D085C085B085A085908580857085608550854085308520851",
			INIT_06 => X"0C700C6F0C6E0C6D0C6C0C6B0C6A0C690C680867086608650864086308620861",
			INIT_07 => X"0C800C7F0C7E0C7D0C7C0C7B0C7A0C790C780C770C760C750C740C730C720C71",
			INIT_08 => X"1090108F108E108D108C108B108A108910881087108610851084108310820C81",
			INIT_09 => X"14A0149F149E149D149C109B109A109910981097109610951094109310921091",
			INIT_0A => X"14B014AF14AE14AD14AC14AB14AA14A914A814A714A614A514A414A314A214A1",
			INIT_0B => X"14C014BF14BE14BD14BC14BB14BA14B914B814B714B614B514B414B314B214B1",
			INIT_0C => X"1CD018CF18CE18CD18CC18CB18CA18C918C818C718C618C518C418C314C214C1",
			INIT_0D => X"1CE01CDF1CDE1CDD1CDC1CDB1CDA1CD91CD81CD71CD61CD51CD41CD31CD21CD1",
			INIT_0E => X"1CF01CEF1CEE1CED1CEC1CEB1CEA1CE91CE81CE71CE61CE51CE41CE31CE21CE1",
			INIT_0F => X"1D001CFF1CFE1CFD1CFC1CFB1CFA1CF91CF81CF71CF61CF51CF41CF31CF21CF1",
			INIT_10 => X"2110210F210E210D210C210B210A2109210821072106210521041D031D021D01",
			INIT_11 => X"2520251F251E251D251C251B251A251925182517251625152114211321122111",
			INIT_12 => X"2930292F292E292D292C292B292A292929282927252625252524252325222521",
			INIT_13 => X"2D402D3F2D3E2D3D2D3C2D3B2D3A2D392D382937293629352934293329322931",
			INIT_14 => X"2D502D4F2D4E2D4D2D4C2D4B2D4A2D492D482D472D462D452D442D432D422D41",
			INIT_15 => X"2D602D5F2D5E2D5D2D5C2D5B2D5A2D592D582D572D562D552D542D532D522D51",
			INIT_16 => X"3570356F356E356D356C356B356A3569396831672D662D652D642D632D622D61",
			INIT_17 => X"3580357F357E357D357C357B357A357935783577357635753574357335723571",
			INIT_18 => X"3590358F358E358D358C358B358A358935883587358635853584358335823581",
			INIT_19 => X"35A0359F359E359D359C359B359A359935983597359635953594359335923591",
			INIT_1A => X"31673167316700003DAC35AB35AA35A935A835A735A635A535A435A335A235A1",
			INIT_1B => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_1C => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_1D => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_1E => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_1F => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_20 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_21 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_22 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_23 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_24 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_25 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_26 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_27 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_28 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_29 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_2A => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_2B => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_2C => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_2D => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_2E => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_2F => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_30 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_31 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_32 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_33 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_34 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_35 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_36 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_37 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_38 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_39 => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_3A => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_3B => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_3C => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_3D => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_3E => X"3167316731673167316731673167316731673167316731673167316731673167",
			INIT_3F => X"3167316731673167316731673167316731673167316731673167316731673167"
		)
-- translate_on
