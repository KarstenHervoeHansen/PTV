-- upconvert.vhd
--
-- Written by:  George Cosens
--              Chief Engineer 
--              Linear Systems Ltd.
--
-- Copyright (c) 2004 Linear Systems Ltd.
-- All rights reserved.
-- Date:  September 29, 2004
--
--
-- This code is intended for use with the Cypress HOTLink II Video Demostration Board
-------------------------------------------------------------------------------------
--
-- This module converts SDI input to HD-SDI output
-- 1080i at 29.97 frames/sec is supported on output for NTSC 270 Mbit/s input
-- clk27 must be syncronous with data_in, clk74 must be derived from clk27 using PLL's
-- for clk27 = 27MHz, clk74 = 74.25/1.001 MHz
--
-- Incoming SDI data is stored in up to 7 line buffers.
-- HDSDI line data is generated by repeating each pixel sample pair twice as follows: 
--   CRnYnCBnYn+1 -> CRnY2nCBnYn+1 CRn+1Yn+1CBn+1Yn+1
-- Lines are repeated as follows:
--    For each 7 lines of SDI data in, the first 6 lines are repeated twice and the 7th line is repeated 3 times.  
--    This generates 15 lines of HDSDI data for each 7 lines of SDI data in. 
--    This stretches the image vertically by about 7% but matches the average line and frame rates for incoming and outgoing data.
-- Unused active video samples in active outgoing video lines are set to black.  
--    This will result in black bars at the sides of the video image.  
--    Some active video lines at the top and bottom of the HDSDI output are not used, they are also set to black. 
--
-- Clocking:
--
-- In order for the up conversion to work I discovered I needed to use both PLL's in the FPGA(U2) connected 
-- in series to get the correct frequency for transmitting.
 
-- The RXCLKB+ input pin of the FPGA is connected to the input of the first PLL in the FPGA. 
-- The FPGA connects the output of the first PLL to  FCLKB+ internally. 
-- The jumper wire connects FCLKB+ output pin of the FPGA to the  RXCLKA+ input pin on the FPGA(U2). 
-- R205 is removed in order to disconnect the RXCLKA+ output pin of the 15G403 chip from the RXCLKA+ input pin of the FPGA(U2). 
-- The RXCLKA+ pin on the FPGA is connected to the input of the second PLL in the FPGA. 
-- The output of the second PLL is connected to FCLKA+ in the FPGA and the inverted output of the PLL is connected to the FCLKA- in the FPGA. 
-- Moving the jumpers on JP11 connects the FCLKA outputs of the FPGA to the REFCLKA inputs of the 15G0403. 
-- The first PLL multiplies  RXCLKB+ by 25/13, The second multiples this result by 10/7.  the resulting frequency is 74.25/1.001 MHz
-- the resulting clock circuit looks like this:
-- 
-- 
--               |------|          |------|  FCLKA+   |------|  REFCLKA+       
--               |      |          |      |---------->|      |----------> 
--  RXCLKB+      |      |  FCLKB+  |      |           |      |        
--  ------------>| PLL1 |--------->| PPL2 |  FCLKA-   | JP11 |  REFCLKA-
--               |      |          |      |---------->|      |----------> 
--               |      |          |      |           |      |        
--               |------|          |------|           |------|

LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;
USE work.pack_crc.all;

ENTITY upconvert IS
	PORT(
		clk27, clk74, reset		: IN	STD_LOGIC;
		data_in					: IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		line_count				: IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		sample_count			: IN	STD_LOGIC_VECTOR(10 DOWNTO 0);
		video_type				: IN	STD_LOGIC_VECTOR(2 DOWNTO 0);
		data_out				: out	STD_LOGIC_VECTOR(19 DOWNTO 0)
	);
END upconvert;
ARCHITECTURE a OF upconvert IS

	component line_buff
		PORT
		(
			data		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
			wren		: IN STD_LOGIC  := '1';
			wraddress		: IN STD_LOGIC_VECTOR (13 DOWNTO 0);
			rdaddress		: IN STD_LOGIC_VECTOR (12 DOWNTO 0);
			wrclock		: IN STD_LOGIC ;
			rdclock		: IN STD_LOGIC ;
			wr_aclr		: IN STD_LOGIC  := '0';
			rd_aclr		: IN STD_LOGIC  := '0';
			q		: OUT STD_LOGIC_VECTOR (19 DOWNTO 0)
		);
	end component;
	
	TYPE IN_STATE_TYPE IS (idle, write);
	SIGNAL instate   : IN_STATE_TYPE;
	SIGNAL wraddress : STD_LOGIC_VECTOR(13 DOWNTO 0);
	signal rdaddress : STD_LOGIC_VECTOR(12 DOWNTO 0);
	signal wrdata : STD_LOGIC_VECTOR(9 DOWNTO 0);
	signal q_sig : STD_LOGIC_VECTOR(19 DOWNTO 0);
	signal bufnum : std_logic_vector(2 downto 0);
	signal wren_sig,ready : STD_LOGIC;

	-- smpte 292 signals
	signal Y_data_out, C_data_out : std_logic_vector(9 downto 0);
	signal linecount : std_logic_vector(10 downto 0);
	signal samplecount, tsamplecount : std_logic_vector(11 downto 0);
	signal xyz : std_logic_vector(9 downto 0);
	signal F,V,H : std_logic;
	signal P : std_logic_vector(3 downto 0);
	signal Y_crc, C_crc : std_logic_vector(17 downto 0);
	signal Y_crc0, C_crc0 : std_logic_vector(17 downto 0);

	-- SMPTE 292 Values for 1080i at 30 fps
	CONSTANT TSL :integer :=2200; -- TOTAL SAMPLES PER LINE
	CONSTANT ASL :integer :=1920; -- ACTIVE SAMPLES PER LINE
	CONSTANT LINES : INTEGER := 1125; -- TOTAL LINES PER FRAME
	CONSTANT VBLANK1A : INTEGER := 20; --  END OF FIRST VERTICAL BALNKING INTERVAL IN FIRST FIELD
	CONSTANT VBLANK1B : INTEGER := 561; --  START OF SECOND VERTICAL BALNKING INTERVAL IN FIRST FIELD
	CONSTANT VBLANK2A : INTEGER := 583; --  END OF FIRST VERTICAL BALNKING INTERVAL IN SECOND FIELD
	CONSTANT VBLANK2B : INTEGER := 1124; --  START OF SECOND VERTICAL BALNKING INTERVAL IN SECOND FIELD

	CONSTANT HALFLINES : INTEGER := LINES/2+1; -- LINES IN FIRST FIELD

	signal line15count : integer range 0 to 14;
	signal rbuf : std_logic_vector(2 downto 0);
	signal y0, y2 : std_logic_vector(9 downto 0);

BEGIN
	process
	begin
		wait until clk74 = '1';
		data_out(19 downto 10) <= Y_data_out;
		data_out(9 downto 0) <= C_data_out;
	end process;
	process(clk27, reset)	-- write process
	begin
	if reset = '1' then
		instate <= idle;
		bufnum <= "000";
		ready <= '0';
	elsif clk27'event and clk27 = '1' then
		CASE instate IS
			WHEN idle =>
				if sample_count = 1441 and line_count = 5 then
					instate <= write;
					bufnum <= "000";
					ready <= '0';
				end if;
			WHEN write =>
				if sample_count = 1441 then
					if line_count = 5 or bufnum >= 6 then
						bufnum <= "000";
					else
						bufnum <= bufnum + 1;
					end if;
				end if;
				if sample_count < 1440 then
					wraddress(13 downto 11) <= bufnum;
					wraddress(10 downto 0) <= sample_count;
					wrdata <= data_in;
					wren_sig <= '1';
				else
					wren_sig <= '0';
				end if;
				if ready = '0' and bufnum = 4 then
					ready <= '1';
				elsif (ready = '1' and sample_count = 1442 and line_count = 5 and bufnum /= 0) then
					ready <= '0';
				end if;
		END CASE;
	end if;
	end process;

	Y_crc0 <= crc_0_4_5_18(Y_data_out,Y_crc);
	C_crc0 <= crc_0_4_5_18(C_data_out,C_crc);
	tsamplecount <= samplecount - 240;
	rdaddress(12 downto 10) <= rbuf;
	rdaddress(9 downto 1) <= tsamplecount(10 downto 2);
	rdaddress(0) <= tsamplecount(0); 
	process (ready,clk74) begin -- read address generator
		if ready = '0' then
			samplecount <= conv_std_logic_vector(ASL,12);
			linecount <= conv_std_logic_vector(1,11);
			rbuf <= "000";
			line15count <= 0;
		elsif clk74'event and clk74 = '1' then
			if samplecount = 1921 then
				case line15count is
					when 0 =>
						line15count <= line15count + 1;
					when 1 =>
						line15count <= line15count + 1;
						rbuf <= rbuf + 1;
					when 2 =>
						line15count <= line15count + 1;
					when 3 =>
						line15count <= line15count + 1;
						rbuf <= rbuf + 1;
					when 4 =>
						line15count <= line15count + 1;
					when 5 =>
						line15count <= line15count + 1;
						rbuf <= rbuf + 1;
					when 6 =>
						line15count <= line15count + 1;
					when 7 =>
						line15count <= line15count + 1;
						rbuf <= rbuf + 1;
					when 8 =>
						line15count <= line15count + 1;
					when 9 =>
						line15count <= line15count + 1;
						rbuf <= rbuf + 1;
					when 10 =>
						line15count <= line15count + 1;
					when 11 =>
						line15count <= line15count + 1;
						rbuf <= rbuf + 1;
					when 12 =>
						line15count <= line15count + 1;
					when 13 =>
						line15count <= line15count + 1;
					when others =>
						line15count <= 0;
						rbuf <= "000";
				end case;
			end if;
			if samplecount = 0 and linecount = 1 and line_count /= 9 then
				linecount <= conv_std_logic_vector(1,11);
				samplecount <= conv_std_logic_vector(0,12);
			elsif samplecount < (TSL-1) then
				samplecount <= samplecount+1;
				if samplecount = (ASL-1) then
					if linecount < LINES then
						linecount <= linecount + 1;
					else
						linecount <= conv_std_logic_vector(1,11);
					end if;
				end if;
			else 
				samplecount <= conv_std_logic_vector(0,12);
			end if;
		end if;
	end process;

	process (ready,clk74) begin -- read process
		if ready = '0' then
			Y_data_out <= "0000000000";
			C_data_out <= "0000000000";
			Y_crc <= conv_std_logic_vector(0,18);
			C_crc <= conv_std_logic_vector(0,18);
		elsif clk74'event and clk74='1' then
			if ((samplecount <= (ASL+6)) and (samplecount > 0)) then
				Y_crc <= crc_0_4_5_18(Y_data_out,Y_crc);
				C_crc <= crc_0_4_5_18(C_data_out,C_crc);
			elsif (samplecount = (ASL+7)) then
				Y_crc <= conv_std_logic_vector(0,18);
				C_crc <= conv_std_logic_vector(0,18);
			end if;
			if samplecount = ASL or samplecount=(TSL-4)then
				Y_data_out <= "1111111111";
				C_data_out <= "1111111111";
			elsif ((samplecount = ASL+1) or (samplecount = ASL+2) or (samplecount = TSL-3) or (samplecount = TSL-2)) then
				Y_data_out <= "0000000000";
				C_data_out <= "0000000000";
			elsif samplecount = ASL+3 or samplecount = TSL-1 then
				Y_data_out <= xyz;
				C_data_out <= xyz;
			ELSIF samplecount = ASL+4 then
				-- LN0 here
				Y_data_out(1 downto 0) <= "00";
				Y_data_out(8 downto 2) <= linecount(6 downto 0);
				Y_data_out(9) <= not linecount(6);
				C_data_out(1 downto 0) <= "00";
				C_data_out(8 downto 2) <= linecount(6 downto 0);
				C_data_out(9) <= not linecount(6);
			ELSIF samplecount = ASL+5 then
				-- LN1 here
				Y_data_out(1 downto 0) <= "00";
				Y_data_out(5 downto 2) <= linecount(10 downto 7);
				Y_data_out(8 downto 6) <= "000";
				Y_data_out(9) <= '1';
				C_data_out(1 downto 0) <= "00";
				C_data_out(5 downto 2) <= linecount(10 downto 7);
				C_data_out(8 downto 6) <= "000";
				C_data_out(9) <= '1';
			elsif samplecount = ASL+6 then
			-- add crc0 here
				Y_Data_out(8 downto 0) <= Y_crc0(8 downto 0);
				Y_data_out(9) <= not Y_crc0(8);
				C_Data_out(8 downto 0) <= C_crc0(8 downto 0);
				C_data_out(9) <= not C_crc0(8);
			elsif samplecount = ASL+7 then
			-- add crc1 here
				Y_Data_out(8 downto 0) <= Y_crc(17 downto 9);
				Y_data_out(9) <= not Y_crc(17);
				C_Data_out(8 downto 0) <= C_crc(17 downto 9);
				C_data_out(9) <= not C_crc(17);
			elsif samplecount > ASL+7 then	-- horizontal blanking interval
				Y_data_out <= "0001000000"; -- 0x040
				C_data_out <= "1000000000"; -- 0x200
			elsif (linecount <= VBLANK1A) or ((linecount >= VBLANK1B) and 
					(linecount <= VBLANK2A)) or (linecount >= VBLANK2B) then -- vertical blanking interval
				Y_data_out <= "0001000000"; -- 0x040
				C_data_out <= "1000000000"; -- 0x200
			else -- active video field
				if samplecount >= 244 and samplecount  < 1680 and 
						((linecount > 37 and linecount < 556) or (linecount > 602 and linecount < 1117) ) then
					Y_data_out <= q_sig(19 downto 10);
					C_data_out <= q_sig(9 downto 0);
				else
					Y_data_out <= conv_std_logic_vector(64,10);--(511,10); --  Y
					C_data_out <= conv_std_logic_vector(512,10);--(512,10); --  Cb or Cr
				end if;
			end if;
		end if;
	end process;

	process (ready,clk74) begin
		if ready = '0' then
			V <= '1';
			F <= '1';
		elsif clk74'event and clk74 = '1' then
			if (linecount <= VBLANK1A) or ((linecount >= VBLANK1B) and (linecount <= VBLANK2A)) or 
					(linecount >= VBLANK2B) then -- vertical blanking interval
				V <= '1';
			else
				V <= '0';
			end if;

			if linecount <= HALFLINES then
				F <= '0';
			else
				F <= '1';
			end if;

			if samplecount > ASL+3 then 
				H <= '0';
			else
				H <= '1';
			end if;
		end if;
	end process;


	xyz(9) <= '1';
	xyz(8) <= F;
	xyz(7) <= V;
	xyz(6) <= H;
	xyz(5 downto 2) <= P;
	xyz(1 downto 0) <= "00";
	WITH xyz(8 downto 6) SELECT
	    p <=
		"0000" WHEN "000",
		"1101" WHEN "001",
		"1011" WHEN "010",
		"0110" WHEN "011",
		"0111" WHEN "100",
		"1010" WHEN "101",
		"1100" WHEN "110",
		"0001" WHEN OTHERS;

	line_buff_inst : line_buff PORT MAP (
			data	 => wrdata,
			wren	 => wren_sig,
			wraddress	 => wraddress,
			rdaddress	 => rdaddress,
			wrclock	 => clk27,
			rdclock	 => clk74,
			wr_aclr	 => reset,
			rd_aclr	 => reset,
			q	 => q_sig
		);

END a;



