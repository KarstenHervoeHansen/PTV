--
-- VROM initialization values for synthesis
-- Created from file NTSC_EG1_RP178.txt on Wed 28 Nov 2001 16:12
-- Formatted for Xilinx XST synthesis tool.
--
attribute WRITE_MODE_A of VROM : label is "READ_FIRST";
attribute WRITE_MODE_B of VROM : label is "READ_FIRST";
attribute INIT_A of VROM : label is "2320D";
attribute INIT_B of VROM : label is "2320D";
attribute SRVAL_A of VROM : label is "2320D";
attribute SRVAL_B of VROM : label is "2320D";
attribute INITP_00 of VROM : label is "000000000000000000000000000000000000000000000000000000155555557E";
attribute INITP_01 of VROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_02 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAFFFFFFFFD4000";
attribute INITP_03 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_04 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAEAAAAAA";
attribute INITP_05 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_06 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_07 of VROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INIT_00 of VROM : label is "0410040F040E040D040C040B040A04090408040704060405040400030002320D";
attribute INIT_01 of VROM : label is "0C200C1F0C1E0C1D0C1C0C1B0C1A0C190C180C170C160C150814041304120411";
attribute INIT_02 of VROM : label is "0C300C2F0C2E0C2D0C2C0C2B0C2A0C290C280C270C260C250C240C230C220C21";
attribute INIT_03 of VROM : label is "0C400C3F0C3E0C3D0C3C0C3B0C3A0C390C380C370C360C350C340C330C320C31";
attribute INIT_04 of VROM : label is "0C500C4F0C4E0C4D0C4C0C4B0C4A0C490C480C470C460C450C440C430C420C41";
attribute INIT_05 of VROM : label is "0C600C5F0C5E0C5D0C5C0C5B0C5A0C590C580C570C560C550C540C530C520C51";
attribute INIT_06 of VROM : label is "0C700C6F0C6E0C6D0C6C0C6B0C6A0C690C680C670C660C650C640C630C620C61";
attribute INIT_07 of VROM : label is "0C800C7F0C7E0C7D0C7C0C7B0C7A0C790C780C770C760C750C740C730C720C71";
attribute INIT_08 of VROM : label is "1090108F108E0C8D0C8C0C8B0C8A0C890C880C870C860C850C840C830C820C81";
attribute INIT_09 of VROM : label is "10A0109F109E109D109C109B109A109910981097109610951094109310921091";
attribute INIT_0A of VROM : label is "10B010AF10AE10AD10AC10AB10AA10A910A810A710A610A510A410A310A210A1";
attribute INIT_0B of VROM : label is "14C014BF14BE14BD14BC14BB14BA14B914B814B710B610B510B410B310B210B1";
attribute INIT_0C of VROM : label is "18D018CF18CE18CD18CC18CB14CA14C914C814C714C614C514C414C314C214C1";
attribute INIT_0D of VROM : label is "18E018DF18DE18DD18DC18DB18DA18D918D818D718D618D518D418D318D218D1";
attribute INIT_0E of VROM : label is "18F018EF18EE18ED18EC18EB18EA18E918E818E718E618E518E418E318E218E1";
attribute INIT_0F of VROM : label is "190018FF18FE18FD18FC18FB18FA18F918F818F718F618F518F418F318F218F1";
attribute INIT_10 of VROM : label is "2110210F210E210D210C210B210A1D091D081907190619051904190319021901";
attribute INIT_11 of VROM : label is "2520251F251E251D251C251B211A211921182117211621152114211321122111";
attribute INIT_12 of VROM : label is "2530252F252E252D252C252B252A252925282527252625252524252325222521";
attribute INIT_13 of VROM : label is "2540253F253E253D253C253B253A253925382537253625352534253325322531";
attribute INIT_14 of VROM : label is "2550254F254E254D254C254B254A254925482547254625452544254325422541";
attribute INIT_15 of VROM : label is "2560255F255E255D255C255B255A255925582557255625552554255325522551";
attribute INIT_16 of VROM : label is "2570256F256E256D256C256B256A256925682567256625652564256325622561";
attribute INIT_17 of VROM : label is "2580257F257E257D257C257B257A257925782577257625752574257325722571";
attribute INIT_18 of VROM : label is "2590258F258E258D258C258B258A258925882587258625852584258325822581";
attribute INIT_19 of VROM : label is "29A0299F299E299D299C299B299A299929982997299629952994299325922591";
attribute INIT_1A of VROM : label is "29B029AF29AE29AD29AC29AB29AA29A929A829A729A629A529A429A329A229A1";
attribute INIT_1B of VROM : label is "2DC02DBF2DBE29BD29BC29BB29BA29B929B829B729B629B529B429B329B229B1";
attribute INIT_1C of VROM : label is "2DD02DCF2DCE2DCD2DCC2DCB2DCA2DC92DC82DC72DC62DC52DC42DC32DC22DC1";
attribute INIT_1D of VROM : label is "31E031DF31DE31DD31DC31DB31DA31D931D831D731D631D531D431D331D231D1";
attribute INIT_1E of VROM : label is "31F031EF31EE31ED31EC31EB31EA31E931E831E731E631E531E431E331E231E1";
attribute INIT_1F of VROM : label is "320031FF31FE31FD31FC31FB31FA31F931F831F731F631F531F431F331F231F1";
attribute INIT_20 of VROM : label is "320D320D0001320D320C320B320A320932083207320632053204320332023201";
attribute INIT_21 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_22 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_23 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_24 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_25 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_26 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_27 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_28 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_29 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_2A of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_2B of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_2C of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_2D of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_2E of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_2F of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_30 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_31 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_32 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_33 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_34 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_35 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_36 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_37 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_38 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_39 of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_3A of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_3B of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_3C of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_3D of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_3E of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
attribute INIT_3F of VROM : label is "320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D";
