		--
		-- Initialize VROM for simulation
		-- Created from file NTSC_EG1_RP178.txt on Wed 28 Nov 2001 16:12
		-- Number of patterns = 2, number of hregion bits = 4, number of vregion bits = 4
		--
-- translate_off
		generic map (
			WRITE_MODE_A => "READ_FIRST",
			WRITE_MODE_B => "READ_FIRST",
			INIT_A       => X"2320D",
			INIT_B       => X"2320D",
			SRVAL_A      => X"2320D",
			SRVAL_B      => X"2320D",
			INITP_00 => X"000000000000000000000000000000000000000000000000000000155555557E",
			INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_02 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAFFFFFFFFD4000",
			INITP_03 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_04 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAEAAAAAA",
			INITP_05 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_06 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INITP_07 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
			INIT_00 => X"0410040F040E040D040C040B040A04090408040704060405040400030002320D",
			INIT_01 => X"0C200C1F0C1E0C1D0C1C0C1B0C1A0C190C180C170C160C150814041304120411",
			INIT_02 => X"0C300C2F0C2E0C2D0C2C0C2B0C2A0C290C280C270C260C250C240C230C220C21",
			INIT_03 => X"0C400C3F0C3E0C3D0C3C0C3B0C3A0C390C380C370C360C350C340C330C320C31",
			INIT_04 => X"0C500C4F0C4E0C4D0C4C0C4B0C4A0C490C480C470C460C450C440C430C420C41",
			INIT_05 => X"0C600C5F0C5E0C5D0C5C0C5B0C5A0C590C580C570C560C550C540C530C520C51",
			INIT_06 => X"0C700C6F0C6E0C6D0C6C0C6B0C6A0C690C680C670C660C650C640C630C620C61",
			INIT_07 => X"0C800C7F0C7E0C7D0C7C0C7B0C7A0C790C780C770C760C750C740C730C720C71",
			INIT_08 => X"1090108F108E0C8D0C8C0C8B0C8A0C890C880C870C860C850C840C830C820C81",
			INIT_09 => X"10A0109F109E109D109C109B109A109910981097109610951094109310921091",
			INIT_0A => X"10B010AF10AE10AD10AC10AB10AA10A910A810A710A610A510A410A310A210A1",
			INIT_0B => X"14C014BF14BE14BD14BC14BB14BA14B914B814B710B610B510B410B310B210B1",
			INIT_0C => X"18D018CF18CE18CD18CC18CB14CA14C914C814C714C614C514C414C314C214C1",
			INIT_0D => X"18E018DF18DE18DD18DC18DB18DA18D918D818D718D618D518D418D318D218D1",
			INIT_0E => X"18F018EF18EE18ED18EC18EB18EA18E918E818E718E618E518E418E318E218E1",
			INIT_0F => X"190018FF18FE18FD18FC18FB18FA18F918F818F718F618F518F418F318F218F1",
			INIT_10 => X"2110210F210E210D210C210B210A1D091D081907190619051904190319021901",
			INIT_11 => X"2520251F251E251D251C251B211A211921182117211621152114211321122111",
			INIT_12 => X"2530252F252E252D252C252B252A252925282527252625252524252325222521",
			INIT_13 => X"2540253F253E253D253C253B253A253925382537253625352534253325322531",
			INIT_14 => X"2550254F254E254D254C254B254A254925482547254625452544254325422541",
			INIT_15 => X"2560255F255E255D255C255B255A255925582557255625552554255325522551",
			INIT_16 => X"2570256F256E256D256C256B256A256925682567256625652564256325622561",
			INIT_17 => X"2580257F257E257D257C257B257A257925782577257625752574257325722571",
			INIT_18 => X"2590258F258E258D258C258B258A258925882587258625852584258325822581",
			INIT_19 => X"29A0299F299E299D299C299B299A299929982997299629952994299325922591",
			INIT_1A => X"29B029AF29AE29AD29AC29AB29AA29A929A829A729A629A529A429A329A229A1",
			INIT_1B => X"2DC02DBF2DBE29BD29BC29BB29BA29B929B829B729B629B529B429B329B229B1",
			INIT_1C => X"2DD02DCF2DCE2DCD2DCC2DCB2DCA2DC92DC82DC72DC62DC52DC42DC32DC22DC1",
			INIT_1D => X"31E031DF31DE31DD31DC31DB31DA31D931D831D731D631D531D431D331D231D1",
			INIT_1E => X"31F031EF31EE31ED31EC31EB31EA31E931E831E731E631E531E431E331E231E1",
			INIT_1F => X"320031FF31FE31FD31FC31FB31FA31F931F831F731F631F531F431F331F231F1",
			INIT_20 => X"320D320D0001320D320C320B320A320932083207320632053204320332023201",
			INIT_21 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_22 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_23 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_24 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_25 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_26 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_27 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_28 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_29 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_2A => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_2B => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_2C => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_2D => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_2E => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_2F => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_30 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_31 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_32 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_33 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_34 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_35 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_36 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_37 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_38 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_39 => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_3A => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_3B => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_3C => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_3D => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_3E => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D",
			INIT_3F => X"320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D320D"
		)
-- translate_on
