--
-- HROM initialization values for synthesis
-- Created from file PAL_EG1_RP178.txt on Fri 27 Aug 2004 14:54
-- Formatted for Xilinx XST synthesis tool.
--
attribute WRITE_MODE_A : string;
attribute WRITE_MODE_B : string;
attribute INIT_A : string;
attribute INIT_B : string;
attribute SRVAL_A : string;
attribute SRVAL_B : string;
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
attribute INIT_00 : string;
attribute INIT_01 : string;
attribute INIT_02 : string;
attribute INIT_03 : string;
attribute INIT_04 : string;
attribute INIT_05 : string;
attribute INIT_06 : string;
attribute INIT_07 : string;
attribute INIT_08 : string;
attribute INIT_09 : string;
attribute INIT_0A : string;
attribute INIT_0B : string;
attribute INIT_0C : string;
attribute INIT_0D : string;
attribute INIT_0E : string;
attribute INIT_0F : string;
attribute INIT_10 : string;
attribute INIT_11 : string;
attribute INIT_12 : string;
attribute INIT_13 : string;
attribute INIT_14 : string;
attribute INIT_15 : string;
attribute INIT_16 : string;
attribute INIT_17 : string;
attribute INIT_18 : string;
attribute INIT_19 : string;
attribute INIT_1A : string;
attribute INIT_1B : string;
attribute INIT_1C : string;
attribute INIT_1D : string;
attribute INIT_1E : string;
attribute INIT_1F : string;
attribute INIT_20 : string;
attribute INIT_21 : string;
attribute INIT_22 : string;
attribute INIT_23 : string;
attribute INIT_24 : string;
attribute INIT_25 : string;
attribute INIT_26 : string;
attribute INIT_27 : string;
attribute INIT_28 : string;
attribute INIT_29 : string;
attribute INIT_2A : string;
attribute INIT_2B : string;
attribute INIT_2C : string;
attribute INIT_2D : string;
attribute INIT_2E : string;
attribute INIT_2F : string;
attribute INIT_30 : string;
attribute INIT_31 : string;
attribute INIT_32 : string;
attribute INIT_33 : string;
attribute INIT_34 : string;
attribute INIT_35 : string;
attribute INIT_36 : string;
attribute INIT_37 : string;
attribute INIT_38 : string;
attribute INIT_39 : string;
attribute INIT_3A : string;
attribute INIT_3B : string;
attribute INIT_3C : string;
attribute INIT_3D : string;
attribute INIT_3E : string;
attribute INIT_3F : string;
attribute WRITE_MODE_A of HROM : label is "READ_FIRST";
attribute WRITE_MODE_B of HROM : label is "READ_FIRST";
attribute INIT_A of HROM : label is "23167";
attribute INIT_B of HROM : label is "23167";
attribute SRVAL_A of HROM : label is "23167";
attribute SRVAL_B of HROM : label is "23167";
attribute INITP_00 of HROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_01 of HROM : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_02 of HROM : label is "5555555555556000000000000000000000000000000000000000000000000000";
attribute INITP_03 of HROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA155555555555555555555555";
attribute INITP_04 of HROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_05 of HROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_06 of HROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INITP_07 of HROM : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
attribute INIT_00 of HROM : label is "0010000F000E000D000C000B000A000900080007000600050004000300020001";
attribute INIT_01 of HROM : label is "0020001F001E001D001C001B001A001900180017001600150014001300120011";
attribute INIT_02 of HROM : label is "0030002F002E002D002C002B002A002900280027002600250024002300220021";
attribute INIT_03 of HROM : label is "0440043F043E043D043C043B043A043904380437043604350434003300320031";
attribute INIT_04 of HROM : label is "0850084F084E084D084C084B084A084908480847084608450844084308420841";
attribute INIT_05 of HROM : label is "0860085F085E085D085C085B085A085908580857085608550854085308520851";
attribute INIT_06 of HROM : label is "0C700C6F0C6E0C6D0C6C0C6B0C6A0C690C680867086608650864086308620861";
attribute INIT_07 of HROM : label is "0C800C7F0C7E0C7D0C7C0C7B0C7A0C790C780C770C760C750C740C730C720C71";
attribute INIT_08 of HROM : label is "1090108F108E108D108C108B108A108910881087108610851084108310820C81";
attribute INIT_09 of HROM : label is "14A0149F149E149D149C109B109A109910981097109610951094109310921091";
attribute INIT_0A of HROM : label is "14B014AF14AE14AD14AC14AB14AA14A914A814A714A614A514A414A314A214A1";
attribute INIT_0B of HROM : label is "14C014BF14BE14BD14BC14BB14BA14B914B814B714B614B514B414B314B214B1";
attribute INIT_0C of HROM : label is "1CD018CF18CE18CD18CC18CB18CA18C918C818C718C618C518C418C314C214C1";
attribute INIT_0D of HROM : label is "1CE01CDF1CDE1CDD1CDC1CDB1CDA1CD91CD81CD71CD61CD51CD41CD31CD21CD1";
attribute INIT_0E of HROM : label is "1CF01CEF1CEE1CED1CEC1CEB1CEA1CE91CE81CE71CE61CE51CE41CE31CE21CE1";
attribute INIT_0F of HROM : label is "1D001CFF1CFE1CFD1CFC1CFB1CFA1CF91CF81CF71CF61CF51CF41CF31CF21CF1";
attribute INIT_10 of HROM : label is "2110210F210E210D210C210B210A2109210821072106210521041D031D021D01";
attribute INIT_11 of HROM : label is "2520251F251E251D251C251B251A251925182517251625152114211321122111";
attribute INIT_12 of HROM : label is "2930292F292E292D292C292B292A292929282927252625252524252325222521";
attribute INIT_13 of HROM : label is "2D402D3F2D3E2D3D2D3C2D3B2D3A2D392D382937293629352934293329322931";
attribute INIT_14 of HROM : label is "2D502D4F2D4E2D4D2D4C2D4B2D4A2D492D482D472D462D452D442D432D422D41";
attribute INIT_15 of HROM : label is "2D602D5F2D5E2D5D2D5C2D5B2D5A2D592D582D572D562D552D542D532D522D51";
attribute INIT_16 of HROM : label is "3570356F356E356D356C356B356A3569396831672D662D652D642D632D622D61";
attribute INIT_17 of HROM : label is "3580357F357E357D357C357B357A357935783577357635753574357335723571";
attribute INIT_18 of HROM : label is "3590358F358E358D358C358B358A358935883587358635853584358335823581";
attribute INIT_19 of HROM : label is "35A0359F359E359D359C359B359A359935983597359635953594359335923591";
attribute INIT_1A of HROM : label is "00003DAF35AE35AD35AC35AB35AA35A935A835A735A635A535A435A335A235A1";
attribute INIT_1B of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_1C of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_1D of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_1E of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_1F of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_20 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_21 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_22 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_23 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_24 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_25 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_26 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_27 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_28 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_29 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_2A of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_2B of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_2C of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_2D of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_2E of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_2F of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_30 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_31 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_32 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_33 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_34 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_35 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_36 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_37 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_38 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_39 of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_3A of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_3B of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_3C of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_3D of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_3E of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
attribute INIT_3F of HROM : label is "3167316731673167316731673167316731673167316731673167316731673167";
