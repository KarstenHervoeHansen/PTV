* C:\PT-Trilevel\pspice\Output-amp.sch

* Schematics Version 9.1 - Web Update 1
* Wed Nov 19 10:19:13 2003



** Analysis setup **
.ac DEC 1000 10 10000K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Output-amp.net"
.INC "Output-amp.als"


.probe


.END
