		--
		-- Initialize CROM for simulation
		-- Created from file PAL_EG1_RP178.txt on Fri 27 Aug 2004 14:54
		-- Number of patterns = 2, number of hregion bits = 4, number of vregion bits = 4
		--
-- translate_off
		generic map (
			WRITE_MODE_A => "READ_FIRST",
			WRITE_MODE_B => "READ_FIRST",
			INIT_A       => X"000",
			INIT_B       => X"000",
			SRVAL_A      => X"000",
			SRVAL_B      => X"000",
			INITP_00 => X"995114445AABBEEF995114445AABBEEF99555555555555559955555555555555",
			INITP_01 => X"995114445AABBEEF995555555555FF11995FF555B5555551995114445AABBEEF",
			INITP_02 => X"0000000000000000995555555555FF11995FF555B5555551995114445AABBEEF",
			INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_04 => X"9955555555555555995555555555555599555555555555559955555555555555",
			INITP_05 => X"9955555555555555995555555555555599555555555555559955555555555555",
			INITP_06 => X"0000000000000000995555555555555599555555555555559955555555555555",
			INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_00 => X"2000200020002000200020002000200020002000200020002000200020002000",
			INIT_01 => X"560000FF6C0000FF200020002000200020002000200020002000200020002000",
			INIT_02 => X"2000200020002000200020002000200020002000200020002000200020002000",
			INIT_03 => X"D80000FFE20000FF200020002000200020002000200020002000200020002000",
			INIT_04 => X"7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800",
			INIT_05 => X"000000FF3A0000FF2000200037F037A837F037A866A866D966A866D966A866D9",
			INIT_06 => X"7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800",
			INIT_07 => X"000000FF3A0000FF2000200037F037A837F037A866A866D966A866D966A866D9",
			INIT_08 => X"7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800",
			INIT_09 => X"000000FF3A0000FF2000200037F037A837F037A866A866D966A866D966A866D9",
			INIT_0A => X"2258222620002000200020007D987D817D987D81200020002000200037F037A8",
			INIT_0B => X"000000FF3A0000FF200020006800680068006800200020002000200020002000",
			INIT_0C => X"2000200020002000462F465C462F465CD600D600D600D6007AC57A327AC57A32",
			INIT_0D => X"000000FF3A0000FF20002000200020002000200031003100200020000E000E00",
			INIT_0E => X"7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800",
			INIT_0F => X"8E0000FFB40000FF2000200037F037A837F037A866A866D966A866D966A866D9",
			INIT_10 => X"7D987D810B670B7E0B670B7E2258222622582226510F5158510F515868006800",
			INIT_11 => X"8E0000FFB40000FF2000200037F037A837F037A866A866D966A866D966A866D9",
			INIT_12 => X"2258222620002000200020007D987D817D987D81200020002000200037F037A8",
			INIT_13 => X"8E0000FFB40000FF200020006800680068006800200020002000200020002000",
			INIT_14 => X"2000200020002000462F465C462F465CD600D600D600D6007AC57A327AC57A32",
			INIT_15 => X"8E0000FFB40000FF20002000200020002000200031003100200020000E000E00",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"2000200020002000200020002000200020002000200020002000200020002000",
			INIT_21 => X"560000FF6C0000FF200020002000200020002000200020002000200020002000",
			INIT_22 => X"2000200020002000200020002000200020002000200020002000200020002000",
			INIT_23 => X"D80000FFE20000FF200020002000200020002000200020002000200020002000",
			INIT_24 => X"CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80",
			INIT_25 => X"000000FF3A0000FF200020004080CC80CC80CC80CC80CC80CC80CC80CC80CC80",
			INIT_26 => X"CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80",
			INIT_27 => X"000000FF3A0000FF20002000CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80",
			INIT_28 => X"8800880088008800880088008800880088008800880088008800880088008800",
			INIT_29 => X"000000FF3A0000FF200020008800880088008800880088008800880088008800",
			INIT_2A => X"8800880088008800880088008800880088008800880088008800880088008800",
			INIT_2B => X"000000FF3A0000FF200020008800880088008800880088008800880088008800",
			INIT_2C => X"8800880088008800880088008800880088008800880088008800880088008800",
			INIT_2D => X"000000FF3A0000FF200020008800880088008800880088008800880088008800",
			INIT_2E => X"CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80",
			INIT_2F => X"8E0000FFB40000FF20002000CC80CC80CC80CC80CC80CC80CC80CC80CC80CC80",
			INIT_30 => X"8800880088008800880088008800880088008800880088008800880088008800",
			INIT_31 => X"8E0000FFB40000FF200020008800880088008800880088008800880088008800",
			INIT_32 => X"8800880088008800880088008800880088008800880088008800880088008800",
			INIT_33 => X"8E0000FFB40000FF200020008800880088008800880088008800880088008800",
			INIT_34 => X"8800880088008800880088008800880088008800880088008800880088008800",
			INIT_35 => X"8E0000FFB40000FF200020008800880088008800880088008800880088008800",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
		)
-- translate_on
