library verilog;
use verilog.vl_types.all;
entity ddr2 is
    generic(
        TCK_MIN         : integer := 5000;
        TJIT_PER        : integer := 125;
        TJIT_DUTY       : integer := 150;
        TJIT_CC         : integer := 250;
        TERR_2PER       : integer := 175;
        TERR_3PER       : integer := 225;
        TERR_4PER       : integer := 250;
        TERR_5PER       : integer := 250;
        TERR_N1PER      : integer := 350;
        TERR_N2PER      : integer := 450;
        TQHS            : integer := 450;
        TAC             : integer := 600;
        TDS             : integer := 150;
        TDH             : integer := 275;
        TDQSCK          : integer := 500;
        TDQSQ           : integer := 350;
        TWPRE           : real    := 0.250000;
        TIS             : integer := 350;
        TIH             : integer := 475;
        TRC             : integer := 55000;
        TRCD            : integer := 15000;
        TWTR            : integer := 10000;
        TRP             : integer := 15000;
        TXARDS          : integer := 6;
        CL_TIME         : integer := 15000;
        AL_MIN          : integer := 0;
        AL_MAX          : integer := 5;
        CL_MIN          : integer := 3;
        CL_MAX          : integer := 6;
        WR_MIN          : integer := 2;
        WR_MAX          : integer := 6;
        BL_MIN          : integer := 4;
        BL_MAX          : integer := 8;
        TCK_MAX         : integer := 8000;
        TCH_MIN         : real    := 0.480000;
        TCH_MAX         : real    := 0.520000;
        TCL_MIN         : real    := 0.480000;
        TCL_MAX         : real    := 0.520000;
        TDIPW           : real    := 0.350000;
        TDQSH           : real    := 0.350000;
        TDQSL           : real    := 0.350000;
        TDSS            : real    := 0.200000;
        TDSH            : real    := 0.200000;
        TWPST           : real    := 0.400000;
        TDQSS           : real    := 0.250000;
        TIPW            : real    := 0.600000;
        TCCD            : integer := 2;
        TRAS_MIN        : integer := 40000;
        TRAS_MAX        : integer := 70000000;
        TRTP            : integer := 7500;
        TWR             : integer := 15000;
        TMRD            : integer := 2;
        TDLLK           : integer := 200;
        TRFC_MIN        : integer := 105000;
        TRFC_MAX        : integer := 70000000;
        TXSRD           : integer := 200;
        TAOND           : integer := 2;
        TAOFD           : real    := 2.500000;
        TAONPD          : integer := 2000;
        TAOFPD          : integer := 2000;
        TANPD           : integer := 3;
        TAXPD           : integer := 8;
        TMOD            : integer := 12000;
        TXARD           : integer := 2;
        TXP             : integer := 2;
        TCKE            : integer := 3;
        DM_BITS         : integer := 2;
        ADDR_BITS       : integer := 13;
        ROW_BITS        : integer := 13;
        COL_BITS        : integer := 10;
        DQ_BITS         : integer := 16;
        DQS_BITS        : integer := 2;
        TRRD            : integer := 10000;
        TFAW            : integer := 50000;
        BA_BITS         : integer := 2;
        MEM_BITS        : integer := 10;
        AP              : integer := 10;
        BL_BITS         : integer := 3;
        BO_BITS         : integer := 2;
        STOP_ON_ERROR   : integer := 1;
        DEBUG           : integer := 1;
        BUS_DELAY       : integer := 0;
        RANDOM_OUT_DELAY: integer := 0;
        RANDOM_SEED     : integer := 711689044;
        RDQSEN_PRE      : integer := 2;
        RDQSEN_PST      : integer := 1;
        RDQS_PRE        : integer := 2;
        RDQS_PST        : integer := 1;
        RDQEN_PRE       : integer := 0;
        RDQEN_PST       : integer := 0;
        WDQS_PRE        : integer := 1;
        WDQS_PST        : integer := 1;
        LOAD_MODE       : integer := 0;
        REFRESH         : integer := 1;
        PRECHARGE       : integer := 2;
        ACTIVATE        : integer := 3;
        WRITE           : integer := 4;
        READ            : integer := 5;
        NOP             : integer := 7;
        PWR_DOWN        : integer := 8;
        SELF_REF        : integer := 9
    );
    port(
        ck              : in     vl_logic;
        ck_n            : in     vl_logic;
        cke             : in     vl_logic;
        cs_n            : in     vl_logic;
        ras_n           : in     vl_logic;
        cas_n           : in     vl_logic;
        we_n            : in     vl_logic;
        dm_rdqs         : inout  vl_logic_vector;
        ba              : in     vl_logic_vector;
        addr            : in     vl_logic_vector;
        dq              : inout  vl_logic_vector;
        dqs             : inout  vl_logic_vector;
        dqs_n           : inout  vl_logic_vector;
        rdqs_n          : out    vl_logic_vector;
        odt             : in     vl_logic
    );
end ddr2;
