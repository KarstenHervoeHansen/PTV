library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity State_timer is
   Port ( f148 :                in    std_logic;
          counter_load :        in    std_logic; -- saetter 'loadable_down_counter' igang
          cnt_load_value :      in    integer range 0 to 1023; -- signal fra 'counter' komponenten - fastsaetter loftet for loadable_down_counter (afhaengigt af positionen i synk signalet)
          cnt_value :           inout integer range 0 to 1023 -- signal til 'state_machine' komponenten

        );
end State_timer;

architecture Behavioral of state_timer is

begin

make_count_down : process(f148)
   begin
      if (f148'event and f148 = '1') then -- debug ( cnt_load_value skifter paa highrising )
         if counter_load = '1' then -- gaa igang ved signal fra tilstandsmaskinen
            cnt_value <= cnt_load_value; -- 'load' taelleren
         else
            if cnt_value /= 0 then
                cnt_value <= (cnt_value -1);
            else
                cnt_value <= 1023;
            end if;
         end if;
      end if;
end process;

end Behavioral;
